`ifndef CFG_SVH
`define CFG_SVH

`define DATA_BITS    8
`define INPUT_BITS   `DATA_BITS
`define OUTPUT_BITS  `DATA_BITS

`endif
