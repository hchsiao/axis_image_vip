`ifndef CFG_SVH
`define CFG_SVH

`define SOURCE_BYTES 1
`define SINK_BYTES   1

`endif
